--=============================================================================
--      File Name: 		
--      	
--      Description:
-- 
--      Version: 1.0
--
--      Created: 
--
--      Last Modified: 
--
--      Compiler: ghdl
--
--      Author: Enrico Tolotto
--
--      University of Udine N° 121127
--============================================================================
